module top_module(
    output zero
);//Build a circuit with no inputs and one output that outputs a constant 0
assign zero = 1'b0;
endmodule
