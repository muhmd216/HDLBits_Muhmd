module top_module( input in, output out );
// assign wire from input to output 
assign out = in ;
endmodule