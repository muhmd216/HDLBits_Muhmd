module top_module( input in, output out );
//implement Not Gate
assign out = ~in ;
endmodule
