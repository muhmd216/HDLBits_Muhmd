module top_module( 
    input a, 
    input b, 
    output out );

//implementation od AND Gate
assign out = a&b ;

endmodule